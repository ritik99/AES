`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:03:43 10/11/2017 
// Design Name: 
// Module Name:    Byte_Sub 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Byte_Sub( data, S, clk);
	input clk; 
	input [127:0]data;
	output reg [127:0]S;
	integer k;
	 
	always@(posedge clk)
	begin
	for(k = 0; k < 120; k = k+8)
		begin
		case(data[k +: 8])
			8'h00: S[k +: 8] = 8'h63;
			8'h01: S[k +: 8] = 8'h7c;
			8'h02: S[k +: 8] = 8'h77;
         8'h03: S[k +: 8] = 8'h7b;
			8'h04: S[k +: 8] = 8'hf2;
			8'h05: S[k +: 8] = 8'h6b;
			8'h06: S[k +: 8] = 8'h6f;
			8'h07: S[k +: 8] = 8'hc5;
			8'h08: S[k +: 8] = 8'h30;
			8'h09: S[k +: 8] = 8'h01;
			8'h0a: S[k +: 8] = 8'h67;
			8'h0b: S[k +: 8] = 8'h2b;
			8'h0c: S[k +: 8] = 8'hfe;
			8'h0d: S[k +: 8] = 8'hd7;
			8'h0e : S[k +: 8] = 8'hab; 
         8'h0f : S[k +: 8] = 8'h76;
			8'h10 : S[k +: 8] = 8'hca;
			8'h11 : S[k +: 8] = 8'h82;
			8'h12 : S[k +: 8] = 8'hc9;
  8'h13 : S[k +: 8] = 8'h7d;
  8'h14 : S[k +: 8] = 8'hfa;
  8'h15 : S[k +: 8] = 8'h59;
  8'h16 : S[k +: 8] = 8'h47;
  8'h17 : S[k +: 8] = 8'hf0;
  8'h18 : S[k +: 8] = 8'had;
  8'h19 : S[k +: 8] = 8'hd4;
  8'h1a : S[k +: 8] = 8'ha2;
  8'h1b : S[k +: 8] = 8'haf;
  8'h1c : S[k +: 8] = 8'h9c;
  8'h1d : S[k +: 8] = 8'ha4;
  8'h1e : S[k +: 8] = 8'h72;
  8'h1f : S[k +: 8] = 8'hc0;
  8'h20 : S[k +: 8] = 8'hb7;
  8'h21 : S[k +: 8] = 8'hfd;
  8'h22 : S[k +: 8] = 8'h93;
  8'h23 : S[k +: 8] = 8'h26;
  8'h24 : S[k +: 8] = 8'h36;
  8'h25 : S[k +: 8] = 8'h3f;
  8'h26 : S[k +: 8] = 8'hf7;
  8'h27 : S[k +: 8] = 8'hcc;
  8'h28 : S[k +: 8] = 8'h34;
  8'h29 : S[k +: 8] = 8'ha5;
  8'h2a : S[k +: 8] = 8'he5;
  8'h2b : S[k +: 8] = 8'hf1;
  8'h2c : S[k +: 8] = 8'h71;
  8'h2d : S[k +: 8] = 8'hd8;
  8'h2e : S[k +: 8] = 8'h31;
  8'h2f : S[k +: 8] = 8'h15;
  8'h30 : S[k +: 8] = 8'h04;
  8'h31 : S[k +: 8] = 8'hc7;
  8'h32 : S[k +: 8] = 8'h23;
  8'h33 : S[k +: 8] = 8'hc3;
  8'h34 : S[k +: 8] = 8'h18;
  8'h35 : S[k +: 8] = 8'h96;
  8'h36 : S[k +: 8] = 8'h05;
  8'h37 : S[k +: 8] = 8'h9a;
  8'h38 : S[k +: 8] = 8'h07;
  8'h39 : S[k +: 8] = 8'h12;
  8'h3a : S[k +: 8] = 8'h80;
  8'h3b : S[k +: 8] = 8'he2;
  8'h3c : S[k +: 8] = 8'heb;
  8'h3d : S[k +: 8] = 8'h27;
  8'h3e : S[k +: 8] = 8'hb2;
  8'h3f : S[k +: 8] = 8'h75;
  8'h40 : S[k +: 8] = 8'h09;
  8'h41 : S[k +: 8] = 8'h83;
  8'h42 : S[k +: 8] = 8'h2c;
  8'h43 : S[k +: 8] = 8'h1a;
  8'h44 : S[k +: 8] = 8'h1b;
  8'h45 : S[k +: 8] = 8'h6e;
  8'h46 : S[k +: 8] = 8'h5a;
  8'h47 : S[k +: 8] = 8'ha0;
  8'h48 : S[k +: 8] = 8'h52;
  8'h49 : S[k +: 8] = 8'h3b;
  8'h4a : S[k +: 8] = 8'hd6;
  8'h4b : S[k +: 8] = 8'hb3;
  8'h4c : S[k +: 8] = 8'h29;
  8'h4d : S[k +: 8] = 8'he3;
  8'h4e : S[k +: 8] = 8'h2f;
  8'h4f : S[k +: 8] = 8'h84;
  8'h50 : S[k +: 8] = 8'h53;
  8'h51 : S[k +: 8] = 8'hd1;
  8'h52 : S[k +: 8] = 8'h00;
  8'h53 : S[k +: 8] = 8'hed;
  8'h54 : S[k +: 8] = 8'h20;
  8'h55 : S[k +: 8] = 8'hfc;
  8'h56 : S[k +: 8] = 8'hb1;
  8'h57 : S[k +: 8] = 8'h5b;
  8'h58 : S[k +: 8] = 8'h6a;
  8'h59 : S[k +: 8] = 8'hcb;
  8'h5a : S[k +: 8] = 8'hbe;
  8'h5b : S[k +: 8] = 8'h39;
  8'h5c : S[k +: 8] = 8'h4a;
  8'h5d : S[k +: 8] = 8'h4c;
  8'h5e : S[k +: 8] = 8'h58;
  8'h5f : S[k +: 8] = 8'hcf;
  8'h60 : S[k +: 8] = 8'hd0;
  8'h61 : S[k +: 8] = 8'hef;
  8'h62 : S[k +: 8] = 8'haa;
  8'h63 : S[k +: 8] = 8'hfb;
  8'h64 : S[k +: 8] = 8'h43;
  8'h65 : S[k +: 8] = 8'h4d;
  8'h66 : S[k +: 8] = 8'h33;
  8'h67 : S[k +: 8] = 8'h85;
  8'h68 : S[k +: 8] = 8'h45;
  8'h69 : S[k +: 8] = 8'hf9;
  8'h6a : S[k +: 8] = 8'h02;
  8'h6b : S[k +: 8] = 8'h7f;
  8'h6c : S[k +: 8] = 8'h50;
  8'h6d : S[k +: 8] = 8'h3c;
  8'h6e : S[k +: 8] = 8'h9f;
  8'h6f : S[k +: 8] = 8'ha8;
  8'h70 : S[k +: 8] = 8'h51;
  8'h71 : S[k +: 8] = 8'ha3;
  8'h72 : S[k +: 8] = 8'h40;
  8'h73 : S[k +: 8] = 8'h8f;
  8'h74 : S[k +: 8] = 8'h92;
  8'h75 : S[k +: 8] = 8'h9d;
  8'h76 : S[k +: 8] = 8'h38;
  8'h77 : S[k +: 8] = 8'hf5;
  8'h78 : S[k +: 8] = 8'hbc;
  8'h79 : S[k +: 8] = 8'hb6;
  8'h7a : S[k +: 8] = 8'hda;
  8'h7b : S[k +: 8] = 8'h21;
  8'h7c : S[k +: 8] = 8'h10;
  8'h7d : S[k +: 8] = 8'hff;
  8'h7e : S[k +: 8] = 8'hf3;
  8'h7f : S[k +: 8] = 8'hd2;
  8'h80 : S[k +: 8] = 8'hcd;
  8'h81 : S[k +: 8] = 8'h0c;
  8'h82 : S[k +: 8] = 8'h13;
  8'h83 : S[k +: 8] = 8'hec;
  8'h84 : S[k +: 8] = 8'h5f;
  8'h85 : S[k +: 8] = 8'h97;
  8'h86 : S[k +: 8] = 8'h44;
  8'h87 : S[k +: 8] = 8'h17;
  8'h88 : S[k +: 8] = 8'hc4;
  8'h89 : S[k +: 8] = 8'ha7;
  8'h8a : S[k +: 8] = 8'h7e;
  8'h8b : S[k +: 8] = 8'h3d;
  8'h8c : S[k +: 8] = 8'h64;
  8'h8d : S[k +: 8] = 8'h5d;
  8'h8e : S[k +: 8] = 8'h19;
  8'h8f : S[k +: 8] = 8'h73;
  8'h90 : S[k +: 8] = 8'h60;
  8'h91 : S[k +: 8] = 8'h81;
  8'h92 : S[k +: 8] = 8'h4f;
  8'h93 : S[k +: 8] = 8'hdc;
  8'h94 : S[k +: 8] = 8'h22;
  8'h95 : S[k +: 8] = 8'h2a;
  8'h96 : S[k +: 8] = 8'h90;
  8'h97 : S[k +: 8] = 8'h88;
  8'h98 : S[k +: 8] = 8'h46;
  8'h99 : S[k +: 8] = 8'hee;
  8'h9a : S[k +: 8] = 8'hb8;
  8'h9b : S[k +: 8] = 8'h14;
  8'h9c : S[k +: 8] = 8'hde;
  8'h9d : S[k +: 8] = 8'h5e;
  8'h9e : S[k +: 8] = 8'h0b;
  8'h9f : S[k +: 8] = 8'hdb;
  8'ha0 : S[k +: 8] = 8'he0;
  8'ha1 : S[k +: 8] = 8'h32;
  8'ha2 : S[k +: 8] = 8'h3a;
  8'ha3 : S[k +: 8] = 8'h0a;
  8'ha4 : S[k +: 8] = 8'h49;
			8'ha5 : S[k +: 8] = 8'h06;
			8'ha6 : S[k +: 8] = 8'h24;
			8'ha7 : S[k +: 8] = 8'h5c;
			8'ha8 : S[k +: 8] = 8'hc2;
			8'ha9 : S[k +: 8] = 8'hd3;
			8'haa : S[k +: 8] = 8'hac;
			8'hab : S[k +: 8] = 8'h62;
			8'hac : S[k +: 8] = 8'h91;
			8'had : S[k +: 8] = 8'h95;
			8'hae : S[k +: 8] = 8'he4;
			8'haf : S[k +: 8] = 8'h79;
			8'hb0 : S[k +: 8] = 8'he7;
			8'hb1 : S[k +: 8] = 8'hc8;
			8'hb2 : S[k +: 8] = 8'h37;
			8'hb3 : S[k +: 8] = 8'h6d;
			8'hb4 : S[k +: 8] = 8'h8d;
			8'hb5 : S[k +: 8] = 8'hd5;
			8'hb6 : S[k +: 8] = 8'h4e;
  			8'hb7 : S[k +: 8] = 8'ha9;
			8'hb8 : S[k +: 8] = 8'h6c;
			8'hb9 : S[k +: 8] = 8'h56;
			8'hba : S[k +: 8] = 8'hf4;
			8'hbb : S[k +: 8] = 8'hea;
			8'hbc : S[k +: 8] = 8'h65;
			8'hbd : S[k +: 8] = 8'h7a;
			8'hbe : S[k +: 8] = 8'hae;
			8'hbf : S[k +: 8] = 8'h08;
			8'hc0 : S[k +: 8] = 8'hba;
			8'hc1 : S[k +: 8] = 8'h78;
			8'hc2 : S[k +: 8] = 8'h25;
			8'hc3 : S[k +: 8] = 8'h2e;
			8'hc4 : S[k +: 8] = 8'h1c;
			8'hc5 : S[k +: 8] = 8'ha6;
			8'hc6 : S[k +: 8] = 8'hb4;
			8'hc7 : S[k +: 8] = 8'hc6;
			8'hc8 : S[k +: 8] = 8'he8;
			8'hc9 : S[k +: 8] = 8'hdd;
			8'hca : S[k +: 8] = 8'h74;
			8'hcb : S[k +: 8] = 8'h1f;
			8'hcc : S[k +: 8] = 8'h4b;
			8'hcd : S[k +: 8] = 8'hbd;
			8'hce : S[k +: 8] = 8'h8b;
			8'hcf : S[k +: 8] = 8'h8a;
			8'hd0 : S[k +: 8] = 8'h70;
			8'hd1 : S[k +: 8] = 8'h3e;
			8'hd2 : S[k +: 8] = 8'hb5;
			8'hd3 : S[k +: 8] = 8'h66;
			8'hd4 : S[k +: 8] = 8'h48;
			8'hd5 : S[k +: 8] = 8'h03;
			8'hd6 : S[k +: 8] = 8'hf6;
			8'hd7 : S[k +: 8] = 8'h0e;
			8'hd8 : S[k +: 8] = 8'h61;
			8'hd9 : S[k +: 8] = 8'h35;
			8'hda : S[k +: 8] = 8'h57;
			8'hdb : S[k +: 8] = 8'hb9;
			8'hdc : S[k +: 8] = 8'h86;
			8'hdd : S[k +: 8] = 8'hc1;
			8'hde : S[k +: 8] = 8'h1d;
			8'hdf : S[k +: 8] = 8'h9e;
			8'he0 : S[k +: 8] = 8'he1;
			8'he1 : S[k +: 8] = 8'hf8;
			8'he2 : S[k +: 8] = 8'h98;
			8'he3 : S[k +: 8] = 8'h11;
			8'he4 : S[k +: 8] = 8'h69;
			8'he5 : S[k +: 8] = 8'hd9;
			8'he6 : S[k +: 8] = 8'h8e;
			8'he7 : S[k +: 8] = 8'h94;
			8'he8 : S[k +: 8] = 8'h9b;
			8'he9 : S[k +: 8] = 8'h1e;
			8'hea : S[k +: 8] = 8'h87;
			8'heb : S[k +: 8] = 8'he9;
			8'hec : S[k +: 8] = 8'hce;
			8'hed : S[k +: 8] = 8'h55;
			8'hee : S[k +: 8] = 8'h28;
			8'hef : S[k +: 8] = 8'hdf;
			8'hf0 : S[k +: 8] = 8'h8c;
			8'hf1 : S[k +: 8] = 8'ha1;
			8'hf2 : S[k +: 8] = 8'h89;
			8'hf3 : S[k +: 8] = 8'h0d;
			8'hf4 : S[k +: 8] = 8'hbf;
			8'hf5 : S[k +: 8] = 8'he6;
			8'hf6 : S[k +: 8] = 8'h42;
			8'hf7 : S[k +: 8] = 8'h68;
			8'hf8 : S[k +: 8] = 8'h41;
			8'hf9 : S[k +: 8] = 8'h99;
			8'hfa : S[k +: 8] = 8'h2d;
			8'hfb : S[k +: 8] = 8'h0f;
			8'hfc : S[k +: 8] = 8'hb0;
			8'hfd : S[k +: 8] = 8'h54;
			8'hfe : S[k +: 8] = 8'hbb;
			8'hff : S[k +: 8] = 8'h16;
		endcase
		end
		end

endmodule